
module test_my_regfile;
    reg [3:0] n1;
    wire [15:0] rd1;

    // レジスタファイルのインスタンス化
    my_regfile uut(.n1(n1), .rd1(rd1));

    // 初期設定とテスト
    initial begin
        $monitor("%t: N1=%d, RD1=%d", $time, n1, rd1);

        n1 = 0;   // 初期値
        #10 n1 = 1;   // 10単位時間後に n1 = 1
        #10 n1 = 2;   // 20単位時間後に n1 = 2
        #10 n1 = 3;   // 30単位時間後に n1 = 3
        #10 n1 = 4;   // 40単位時間後に n1 = 4
        #10 n1 = 5;   // 50単位時間後に n1 = 5
        #10 n1 = 6;   // 60単位時間後に n1 = 6
        #10 n1 = 7;   // 70単位時間後に n1 = 7
        #10 n1 = 8;   // 80単位時間後に n1 = 8
        #10 n1 = 9;   // 90単位時間後に n1 = 9
        #10 $finish;  // シミュレーション終了
    end
endmodule
