module my_alu1 ( cin, a, b, r, cout, s_sub, s_fas, s_and, s_or, s_xor, s_not);
input   cin, a, b, s_sub, s_fas, s_and, s_or, s_xor, s_not;
output  r, cout;
wire r_in;

// <<ここを埋めよ. Please fill in here>>

endmodule

